`default_nettype none



module uart_axis (
	input logic in
	output logic out);

	assign out = in;


endmodule
