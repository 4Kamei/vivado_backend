typedef logic [7:0] device_type;
localparam device_type CLOCK_COUNTER_DEVICE_TYPE = 8'h01;   //{"display": "Clock Counter"}
localparam device_type I2C_MASTER_DEVICE_TYPE    = 8'h02;   //{"display": "I2C Master"}
localparam device_type REGISTER_MAP_DEVICE_TYPE  = 8'h03;   //{"display": "Register Map"}
    
