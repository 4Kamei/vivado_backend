localparam logic [7:0] AXIS_DEBUG_IDS_CLK_LOGIC     = 8'h00;
localparam logic [7:0] AXIS_DEBUG_IDS_CLK_QSFP      = 8'h01;
localparam logic [7:0] AXIS_DEBUG_IDS_CLK_GTX_REF   = 8'h02;
localparam logic [7:0] AXIS_DEBUG_IDS_CLK_GTX_TX    = 8'h03;
localparam logic [7:0] AXIS_DEBUG_IDS_CLK_PCS_TX    = 8'h04;
localparam logic [7:0] AXIS_DEBUG_IDS_CLK_FABRIC_TX = 8'h05;
localparam logic [7:0] AXIS_DEBUG_IDS_CLK_GTX_RX    = 8'h06;

//I2C
localparam logic [7:0] AXIS_DEBUG_IDS_I2C_TEMP      = 8'h00;

//Register map
localparam logic [7:0] AXIS_DEBUG_IDS_REGISTER_MAP  = 8'h00;
