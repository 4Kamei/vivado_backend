module IBUFGDS (
        input wire I,
        input wire IB,
        output wire O
    );

    assign O = I;

endmodule
